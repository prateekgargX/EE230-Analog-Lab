Inverting Schimdt trigger B
*Including the predefined op-amp subcircuit file
.include ua741.txt
.include zener_1N4732A.txt
.include Diode_1N914.txt
*Connections as mentioned in subcircuit file
x1 8 2 3 4 5 UA741
vcc 3 0 dc 15v
vee 4 0 dc -15v
R1 3 6 13.3k
R2 4 7 13.3k
D1 6 5 1N914
D2 6 8 1N914
D3 5 7 1N914
D4 8 7 1N914
XZ1 9 8 DI_1N4732A
XZ2 9 0 DI_1N4732A
vin 2 0 dc 0

.dc vin -10 10 0.01
.dc vin 10 -10 -0.01 
.control
run
plot dc2.v(8) dc1.v(8)
*print dc2.v(7) 
*print dc1.v(7)
.endc
.end

