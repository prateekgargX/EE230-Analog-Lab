RC Bandpass Filter
*describe circuit
* <element-name> <nodes> <value/nodel>
r1 1 2 10k
c1 2 3 0.1u
r2 3 0 10k
c2 3 0 0.1u
v 1 0 dc 0 ac 1 $ac analysis
*analysis command
.ac dec 20 0.1u 100Meg 

.control 
run

*display cmd
plot vdb(3)
print vdb(3)
*end control mode
.endc 

*end netlist
.end