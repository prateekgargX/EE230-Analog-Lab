RC Highpass Filter
*describe circuit
* <element-name> <nodes> <value/nodel>
c 1 2 0.1u
r 2 0 10k
v 1 0 dc 0 ac 1 $ac analysis
*analysis command
.ac dec 10 1 10Meg

.control 
run

*display cmd
plot vdb(2)
print vdb(2)  
*end control mode
.endc 

*end netlist
.end