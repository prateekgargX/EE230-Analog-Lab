RLC Bandpass Filter
*describe circuit
* <element-name> <nodes> <value/nodel>
l 1 2 10m
c 2 3 0.1u
r 3 0 1k

v 1 0 dc 0 ac 1 $ac analysis
*analysis command
.ac dec 20 0.1u 100Meg 

.control 
run

*display cmd
plot vdb(3)
print vdb(3)
*end control mode
.endc 

*end netlist
.end