Op-amp 741 based circuit-3
*Including the predefined op-amp subcircuit file
.include ua741.txt
.include zener_B.txt

.SUBCKT ZENER_12 1 2
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 3.48
.MODEL DF D ( IS=27.5p RS=0.620 N=1.10 CJO=78.3p VJ=1.00 M=0.330
+ TT=50.1n)
.MODEL DR D ( IS=5.49f RS=50 N=1.77 )
.ENDS

*Connections as mentioned in subcircuit file
x1 2 0 3 4 5 UA741
R1 2 6 8.2K
R2 2 7 15K 
R3 5 7 1K
xz1 8 7 ZENER_12
xz2 8 0 ZENER_12
vcc 3 0 dc 15v
vee 4 0 dc -15v
* vin 6 0 sin(0 5 1k 0 0)
* .tran 0.0001m 0.01 

* .control
* run
* plot v(7) vs v(6) 
* plot v(7) v(6) 

vin 6 0 dc 0 ac 5

.dc vin -5 5 0.01
.dc vin 5 -5 -0.01 
.control
run
plot dc2.v(7) dc1.v(7)
*print dc2.v(7) 
*print dc1.v(7)
.endc
.end