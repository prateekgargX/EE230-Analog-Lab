RC circuit transient analysis
*tau =1m

*describe circuit
* <element-name> <nodes> <value/nodel>
r 1 2 10k
c 2 0 0.1u
*v 1 0 pwl(0 0 10m 0 10.9999m 0 11m 5 20m 5 20.00001m 0)
v 1 0 pulse(0 5 0 0 0 10m 20m)
*analysis command
.tran 1m 100m 

.control 
run

*display cmd
plot v(1) v(2)
print v(2)
*end control mode
.endc 

*end netlist
.end