Family of Curves
*Model file for the MOSFET
.include tsmc_spice_180nm.txt
*Usually, the order of terminals are
*drain, gate, source and body respectively
m1 d g gnd gnd CMOSN
vgs g gnd dc 1.8V
vds dummy gnd dc 1.8V
vdummy dummy d dc 0V
.control
dc vds 0 1.8 0.02 vgs 0 1 0.2
plot i(vdummy)
.endc
.end