RC Lowpass Filter

*describe circuit
* <element-name> <nodes> <value/nodel>
r 1 2 10k
c 2 0 0.1u
vin 1 0 dc 0 ac 1 $ac analysis
*analysis command
.ac dec 10 1 10Meg 

.control 
run

*display cmd
plot vdb(2)
print vdb(2)
*end control mode
.endc 

*end netlist
.end