Bridge-Rectifier circuit
.include 1N4007.txt

*describe circuit
* <element-name> <nodes> <value/nodel>

d1 1 4 DI_1N4007
vd1 4 3 dc 0

d2 0 1 DI_1N4007
d3 2 5 DI_1N4007
vd3 5 3

d4 0 2 DI_1N4007
r1 3 0 1k

vin 1 2 sin(0 21.21320 50 0 0)

*analysis command
.tran 0.0005 0.2

.control 
run

*display cmd
plot v(3) 
*v(1,2)
plot i(vd1) i(vd3)
print v(3) > voltage
print i(vd1) i(vd3) >current
*end control mode
.endc 

*end netlist
.end