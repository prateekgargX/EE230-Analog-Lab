Op-amp 741 based circuit-4
*Including the predefined op-amp subcircuit file
.include ua741.txt
.include zener_B.txt

.SUBCKT ZENER_12 1 2
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 3.58
.MODEL DF D ( IS=27.5p RS=0.620 N=1.10 CJO=78.3p VJ=1.00 M=0.330
+ TT=50.1n)
.MODEL DR D ( IS=5.49f RS=50 N=1.77 )
.ENDS

.SUBCKT Circuit_1 IN OUT COMM
x1 2 COMM 3 4 5 UA741
R1 2 IN 8.2K
R2 2 OUT 15K 
R3 5 OUT 1K
xz1 8 OUT ZENER_12
xz2 8 COMM ZENER_12
vcc 3 COMM dc 15v
vee 4 COMM dc -15v
.ENDS

.SUBCKT Circuit_2 IN OUT COMM
x1 COMM 2 3 4 OUT UA741
c1 2 OUT 47n
r1 2 OUT 1.5Meg
r2 2 IN 18k
vcc 3 COMM dc 15v
vee 4 COMM dc -15v
.ENDS

x5 1 2 0 Circuit_1
x8 2 1 0 Circuit_2
*vin 1 0 sin(0 5 1k 0 0)
.tran 0.001m 105m 95m
.control
run
plot v(2) v(1)
*print v(2) v(1) 
.endc
.end
