Schmitt trigger
*Including the predefined op-amp subcircuit file
.include ua741.txt
.include zener_B.txt

.SUBCKT ZENER_12 1 2
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 3.48
.MODEL DF D ( IS=27.5p RS=0.620 N=1.10 CJO=78.3p VJ=1.00 M=0.330
+ TT=50.1n)
.MODEL DR D ( IS=5.49f RS=50 N=1.77 )
.ENDS

*Connections as mentioned in subcircuit file
x1 2 9 3 4 5 UA741
R1 2 6 10K
R2 2 7 10K 
R3 5 7 1K
xz1 8 7 ZENER_12
xz2 8 0 ZENER_12
vcc 3 0 dc 15v
vee 4 0 dc -15v

va 6 0 dc 3
vin 9 0 sin(0 6 1k 0 0)
.tran 0.001m 0.01
.control
run
plot v(7) vs v(9)
plot v(7) v(9)
*print v(9) v(7)
.endc
.end