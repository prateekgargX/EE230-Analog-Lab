Inverting-Amplifier using op-amp 741
*Including the predefined op-amp subcircuit file
.include ua741.txt
*Connections as mentioned in subcircuit file
x1 0 1 2 3 4 UA741
r1 5 1 10k
rt 4 1 470k
c1 4 1 0.01u
vcc 2 0 dc 15v
vee 3 0 dc -15v
*Giving a sinusoidal input
*vin 5 0 sin (0 0.1 1k 0 0)
vin 5 0 pulse (2 -2 0 1p 1p 0.5m 1m)
.tran 0.02ms 20ms
.control
run
plot v(5) v(4)
.endc