Opamp lm324 based circuit-1
*Including the predefined op-amp subcircuit file
.include lm324.txt
.include ua741.txt

*Connections as mentioned in subcircuit file
x1 1 2 3 0 4 LM324
*x1 1 2 3 0 4 ua741
rg 2 5 20k
rf 2 4 180k
rl 4 0 10k
r1 6 5 75k
r2 0 5 820
c1 3 0 0.01
c2 0 5 0.01
vr1 6 0 dc 5
vcc 3 0 dc 5
vin 1 0 dc 0
.dc vin 0.1 5 0.1
.control
run
plot v(4) v(1)
*print v(4) v(1)
.endc   
.end